Vim�UnDo� ��@6��p�GbQ�*�Ym��ҳ4}��ݾ�$�      input 	[32:0]	RS2_Data_i;      	                       a�:&    _�                             ����                                                                                                                                                                                                                                                                                                                                                             a���     �                   5��                                                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a���     �                  module Equal();5��                                                �                                                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             a���     �                5��                                                �                                             �                                             �                     	                 	       �                                              �                                               �                     
                 
       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a���     �               	RS1_Data_i5��                                             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a���     �               	RS2_Data_i5��                         &                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a���     �               	�             5��                          (                      �                         )                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a���     �                  �               5��                          3                      �                          3                      �                       	   4               	       5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             a��     �                 	input 	[]5��                         <                      5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             a��	     �                 input 	[31:0]5��                         A                      �                        B                     5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             a��     �                  �               5��                          N                      �                          N                      �                         N                     �                         N                     �                      	   N              	       5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             a��     �                 	input 	[]5��                         V                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��     �               input 	[31:0] RS1_Data_i;5��                         A                      5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��     �               input 	[31:0]	 RS1_Data_i;5��                        A                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��    �                 input 	[32:0]5��                         [                      �                     
   \              
       �              
          \       
              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��    �                  �               5��                          h                      �                       
   h               
       �                        p                     5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                                             a��W     �   	               �   	            5��    	                      x                      �    	                      x                      �    
                   	   y               	       5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                                             a��[     �   
             �   
          5��    
                      y                      �    
                      y                      �    
                    z                     �    
                    �                     5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             a��c     �   
            assign data_o = ()5��    
                     �                      �    
                    �                     �    
                 
   �              
       �    
          
       
   �       
       
       5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                                             a��i     �   
            *assign data_o = (RS1_Data_i == RS2_Data_i)5��    
   *                  �                      5�_�                       6    ����                                                                                                                                                                                                                                                                                                                                                             a��v    �                �             5��                          �                      �                          �                      �                          �                      5�_�                        	    ����                                                                                                                                                                                                                                                                                                                                                             a�:%    �      	         input 	[32:0]	RS2_Data_i;5��       	                 W                     5��